Teensy-Theremin5 -3
R8 8 3 10k
R9 11 3 10k
R7 9 3 10k
R10 10 3 10k
R2 3 13 10k

.TRAN 1ms 100ms
* .AC DEC 100 100 1MEG
.END
